`timescale 1 ns/ 10 ps
module tb_contadorpulsos;
reg push;
wire [7:0] contador2;

localparam periodo = 20;
localparam medioperiodo=periodo/2;

contadorpulsos DUT1(.entrada(push), .contador(contador2) );

always 
	#periodo push=~push;

initial
begin
	$display("***************Iniciando simulacion***************");
	push=0;
	#medioperiodo;
	$monitor($time, "reloj = %b, contador=%d", push, contador2);
end	
endmodule

